//////////////////////////////////////////////////////////////////////////////////
// Company:Meyesemi 
// Engineer: Will
// 
// Create Date: 2023-03-17  
// Design Name:  
// Module Name: 
// Project Name: 
// Target Devices: Pango
// Tool Versions: 
// Description: 
//      
// Dependencies: 
// 
// Revision:
// Revision 1.0 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
//sclk，sdin数据传输时序代码（i2c写控制代码）
module i2c_com (
    input clock_i2c,  //i2c控制接口传输所需时钟，0-400khz，此处为20khz
    input clock_i2c_opposite,  //i2c控制接口传输所需时钟，0-400khz，此处为20khz

    input camera_rstn,
    output ack,  //应答信号
    input [31:0] i2c_data,  //sdin接口传输的32位数据
    input start,  //开始传输标志
    output reg tr_end,  //传输结束标志
    output i2c_sclk,  //FPGA与camera iic时钟接口
    inout i2c_sdat  //FPGA与camera iic数据接口
);

  reg [5:0] cyc_count;
  reg reg_sdat;
  reg sclk;
  reg ack1, ack2, ack3;


  assign ack = ack1 | ack2 | ack3;
  assign i2c_sdat = reg_sdat ? 1'bz : 0;

  assign i2c_sclk = sclk | (((cyc_count >= 4) & (cyc_count <= 39)) ? clock_i2c_opposite : 0);

  // wire ce1, ce2;
  // wire clk_temp;
  // assign ce1 = ((cyc_count >= 4) & (cyc_count <= 39)) ? 1 : 0;
  // assign ce2 = ~sclk;
  // GTP_CLKBUFGCE #(
  //     .DEFAULT_VALUE(1'b0)  //1'b0; 1'b1
  // ) GTP_CLKBUFGCE_SCLK0 (
  //     .CLKIN(clock_i2c_opposite),
  //     .CE(ce1),
  //     .CLKOUT(clk_temp)
  // );

  // GTP_CLKBUFGCE #(
  //     .DEFAULT_VALUE(1'b1)  //1'b0; 1'b1
  // ) GTP_CLKBUFGCE_SCLK1 (
  //     .CLKIN(clk_temp),
  //     .CE(ce2),
  //     .CLKOUT(i2c_sclk)
  // );



  always @(posedge clock_i2c) begin
    if (!camera_rstn) cyc_count <= 6'b111111;
    else begin
      if (start == 0) cyc_count <= 0;
      else if (cyc_count < 6'b111111) cyc_count <= cyc_count + 1;
    end
  end


  always @(posedge clock_i2c) begin
    if (!camera_rstn) begin
      tr_end <= 0;
      ack1 <= 1;
      ack2 <= 1;
      ack3 <= 1;
      sclk <= 1;
      reg_sdat <= 1;
    end else
      case (cyc_count)
        0: begin
          ack1 <= 1;
          ack2 <= 1;
          ack3 <= 1;
          tr_end <= 0;
          sclk <= 1;
          reg_sdat <= 1;
        end
        1:  reg_sdat <= 0;  //开始传输
        2:  sclk <= 0;
        3:  reg_sdat <= i2c_data[31];
        4:  reg_sdat <= i2c_data[30];
        5:  reg_sdat <= i2c_data[29];
        6:  reg_sdat <= i2c_data[28];
        7:  reg_sdat <= i2c_data[27];
        8:  reg_sdat <= i2c_data[26];
        9:  reg_sdat <= i2c_data[25];
        10: reg_sdat <= i2c_data[24];
        11: reg_sdat <= 1;  //应答信号
        12: begin
          reg_sdat <= i2c_data[23];
          ack1 <= i2c_sdat;
        end
        13: reg_sdat <= i2c_data[22];
        14: reg_sdat <= i2c_data[21];
        15: reg_sdat <= i2c_data[20];
        16: reg_sdat <= i2c_data[19];
        17: reg_sdat <= i2c_data[18];
        18: reg_sdat <= i2c_data[17];
        19: reg_sdat <= i2c_data[16];
        20: reg_sdat <= 1;  //应答信号       
        21: begin
          reg_sdat <= i2c_data[15];
          ack1 <= i2c_sdat;
        end
        22: reg_sdat <= i2c_data[14];
        23: reg_sdat <= i2c_data[13];
        24: reg_sdat <= i2c_data[12];
        25: reg_sdat <= i2c_data[11];
        26: reg_sdat <= i2c_data[10];
        27: reg_sdat <= i2c_data[9];
        28: reg_sdat <= i2c_data[8];
        29: reg_sdat <= 1;  //应答信号       
        30: begin
          reg_sdat <= i2c_data[7];
          ack2 <= i2c_sdat;
        end
        31: reg_sdat <= i2c_data[6];
        32: reg_sdat <= i2c_data[5];
        33: reg_sdat <= i2c_data[4];
        34: reg_sdat <= i2c_data[3];
        35: reg_sdat <= i2c_data[2];
        36: reg_sdat <= i2c_data[1];
        37: reg_sdat <= i2c_data[0];
        38: reg_sdat <= 1;  //应答信号       
        39: begin
          ack3 <= i2c_sdat;
          sclk <= 0;
          reg_sdat <= 0;
        end
        40: sclk <= 1;
        41: begin
          reg_sdat <= 1;
          tr_end   <= 1;
        end
      endcase

  end
endmodule
